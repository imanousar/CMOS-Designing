magic
tech scmos
timestamp 1594160246
<< nwell >>
rect 29 -6 312 26
rect 78 -68 104 -6
rect 140 -68 166 -6
rect 209 -68 235 -6
rect 280 -7 312 -6
rect 280 -68 310 -7
<< polysilicon >>
rect 31 4 33 6
rect 38 4 66 6
rect 71 4 127 6
rect 137 4 191 6
rect 211 4 245 6
rect 285 4 312 6
rect 41 -10 43 4
rect 38 -12 43 -10
rect 49 -23 52 -21
rect 62 -23 64 -21
rect 70 -23 80 -21
rect 100 -23 102 -21
rect 111 -23 114 -21
rect 124 -23 126 -21
rect 132 -23 142 -21
rect 162 -23 164 -21
rect 180 -23 184 -21
rect 194 -23 196 -21
rect 202 -23 212 -21
rect 232 -23 234 -21
rect 70 -25 72 -23
rect 132 -25 134 -23
rect 202 -25 204 -23
rect 248 -26 251 -24
rect 261 -26 264 -24
rect 275 -26 284 -24
rect 304 -26 307 -24
rect 275 -29 277 -26
rect 271 -31 277 -29
rect 49 -51 52 -49
rect 62 -51 80 -49
rect 100 -51 102 -49
rect 111 -51 115 -49
rect 125 -51 142 -49
rect 162 -51 164 -49
rect 180 -51 185 -49
rect 195 -51 212 -49
rect 232 -51 234 -49
rect 248 -51 251 -49
rect 261 -51 284 -49
rect 304 -51 307 -49
<< ndiffusion >>
rect 52 -21 62 -19
rect 114 -21 124 -19
rect 184 -21 194 -19
rect 52 -25 62 -23
rect 114 -25 124 -23
rect 184 -25 194 -23
rect 251 -24 261 -22
rect 251 -28 261 -26
rect 52 -49 62 -47
rect 52 -53 62 -51
rect 115 -49 125 -47
rect 115 -53 125 -51
rect 185 -49 195 -47
rect 185 -53 195 -51
rect 251 -49 261 -47
rect 251 -53 261 -51
<< pdiffusion >>
rect 33 6 38 8
rect 66 6 71 8
rect 127 6 137 9
rect 191 6 211 9
rect 245 6 285 10
rect 33 2 38 4
rect 66 2 71 4
rect 127 1 137 4
rect 191 1 211 4
rect 245 2 285 4
rect 80 -21 100 -19
rect 142 -21 162 -19
rect 212 -21 232 -19
rect 80 -25 100 -23
rect 142 -25 162 -23
rect 212 -25 232 -23
rect 284 -24 304 -22
rect 284 -28 304 -26
rect 80 -49 100 -47
rect 80 -52 100 -51
rect 142 -49 162 -47
rect 142 -52 162 -51
rect 212 -49 232 -46
rect 212 -52 232 -51
rect 284 -49 304 -46
rect 284 -52 304 -51
<< metal1 >>
rect 30 18 86 19
rect 30 14 46 18
rect 50 14 57 18
rect 61 14 86 18
rect 30 13 86 14
rect 94 18 149 19
rect 94 14 118 18
rect 122 14 149 18
rect 94 13 149 14
rect 157 18 222 19
rect 157 14 183 18
rect 187 14 222 18
rect 157 13 222 14
rect 229 18 298 19
rect 229 14 234 18
rect 238 14 298 18
rect 229 13 245 14
rect 34 -9 38 -3
rect 34 -16 38 -13
rect 67 -15 71 -3
rect 88 -4 92 13
rect 128 -15 133 -3
rect 151 -4 155 13
rect 223 -3 228 13
rect 285 13 298 14
rect 304 13 312 19
rect 45 -20 49 -16
rect 62 -19 80 -15
rect 107 -19 111 -15
rect 124 -19 142 -15
rect 175 -18 180 -14
rect 198 -15 203 -3
rect 194 -19 212 -15
rect 243 -22 248 -17
rect 265 -18 270 -2
rect 299 -3 303 13
rect 261 -22 284 -18
rect 62 -29 68 -25
rect 124 -29 130 -25
rect 194 -29 200 -25
rect 86 -33 94 -30
rect 151 -33 158 -30
rect 55 -34 94 -33
rect 55 -38 63 -34
rect 67 -38 94 -34
rect 55 -43 58 -38
rect 86 -41 94 -38
rect 119 -37 126 -33
rect 130 -37 158 -33
rect 222 -34 229 -29
rect 261 -32 267 -28
rect 119 -38 158 -37
rect 119 -43 122 -38
rect 151 -42 158 -38
rect 190 -38 196 -34
rect 200 -38 229 -34
rect 294 -36 304 -32
rect 190 -43 193 -38
rect 222 -41 229 -38
rect 254 -40 272 -36
rect 276 -40 304 -36
rect 254 -43 259 -40
rect 284 -41 304 -40
rect 20 -58 25 -53
rect 45 -56 49 -52
rect 55 -68 59 -57
rect 107 -56 111 -52
rect 13 -82 20 -79
rect 55 -79 59 -72
rect 86 -64 94 -58
rect 175 -56 180 -52
rect 86 -68 98 -64
rect 118 -66 122 -57
rect 118 -79 122 -70
rect 149 -63 157 -57
rect 243 -56 248 -52
rect 149 -68 161 -63
rect 188 -65 192 -57
rect 221 -62 229 -57
rect 217 -68 229 -62
rect 188 -79 192 -69
rect 255 -67 259 -57
rect 296 -62 304 -57
rect 291 -68 304 -62
rect 255 -79 259 -71
rect 25 -82 63 -79
rect 67 -82 274 -79
rect 247 -102 284 -98
<< metal2 >>
rect 45 -20 49 -16
rect 20 -77 25 -63
rect 34 -77 38 -20
rect 45 -56 49 -24
rect 45 -68 49 -60
rect 68 -93 72 -25
rect 86 -68 94 13
rect 107 -19 111 -15
rect 107 -56 111 -23
rect 107 -68 111 -60
rect 130 -93 134 -25
rect 149 -68 157 13
rect 175 -56 180 -14
rect 175 -68 180 -60
rect 200 -93 204 -25
rect 222 -68 229 13
rect 243 -56 248 -17
rect 243 -68 248 -60
rect 267 -93 271 -28
rect 298 -68 304 13
rect 68 -98 247 -93
rect 252 -98 284 -93
<< ntransistor >>
rect 52 -23 62 -21
rect 114 -23 124 -21
rect 184 -23 194 -21
rect 251 -26 261 -24
rect 52 -51 62 -49
rect 115 -51 125 -49
rect 185 -51 195 -49
rect 251 -51 261 -49
<< ptransistor >>
rect 33 4 38 6
rect 66 4 71 6
rect 127 4 137 6
rect 191 4 211 6
rect 245 4 285 6
rect 80 -23 100 -21
rect 142 -23 162 -21
rect 212 -23 232 -21
rect 284 -26 304 -24
rect 80 -51 100 -49
rect 142 -51 162 -49
rect 212 -51 232 -49
rect 284 -51 304 -49
<< polycontact >>
rect 34 -13 38 -9
rect 45 -24 49 -20
rect 107 -23 111 -19
rect 175 -23 180 -18
rect 68 -29 72 -25
rect 130 -29 134 -25
rect 200 -29 204 -25
rect 243 -27 248 -22
rect 267 -32 271 -28
rect 45 -52 49 -48
rect 107 -52 111 -48
rect 175 -52 180 -47
rect 243 -52 248 -47
<< ndcontact >>
rect 52 -19 62 -15
rect 114 -19 124 -15
rect 184 -19 194 -15
rect 251 -22 261 -18
rect 52 -29 62 -25
rect 114 -29 124 -25
rect 184 -29 194 -25
rect 251 -32 261 -28
rect 52 -47 62 -43
rect 115 -47 125 -43
rect 52 -57 62 -53
rect 185 -47 195 -43
rect 115 -57 125 -53
rect 251 -47 261 -43
rect 185 -57 195 -53
rect 251 -57 261 -53
<< pdcontact >>
rect 33 8 39 13
rect 66 8 72 13
rect 127 9 137 13
rect 191 9 211 13
rect 245 10 285 14
rect 33 -3 39 2
rect 66 -3 72 2
rect 127 -3 137 1
rect 191 -3 211 1
rect 245 -2 285 2
rect 80 -19 100 -15
rect 142 -19 162 -15
rect 212 -19 232 -15
rect 80 -30 100 -25
rect 142 -30 162 -25
rect 212 -29 232 -25
rect 284 -22 304 -18
rect 284 -32 304 -28
rect 80 -47 100 -41
rect 142 -47 162 -42
rect 80 -58 100 -52
rect 212 -46 232 -41
rect 142 -57 162 -52
rect 284 -46 304 -41
rect 212 -57 232 -52
rect 284 -57 304 -52
<< m2contact >>
rect 86 13 94 19
rect 149 13 157 19
rect 222 13 229 19
rect 34 -20 38 -16
rect 45 -16 49 -12
rect 107 -15 111 -11
rect 298 13 304 19
rect 175 -14 180 -10
rect 243 -17 248 -12
rect 20 -63 25 -58
rect 45 -60 49 -56
rect 20 -82 25 -77
rect 107 -60 111 -56
rect 86 -73 94 -68
rect 175 -60 180 -56
rect 243 -60 248 -56
rect 149 -73 157 -68
rect 222 -74 229 -68
rect 298 -74 304 -68
rect 247 -98 252 -93
<< psubstratepcontact >>
rect 63 -38 67 -34
rect 126 -37 130 -33
rect 196 -38 200 -34
rect 272 -40 276 -36
rect 20 -53 25 -48
rect 55 -72 59 -68
rect 118 -70 122 -66
rect 188 -69 192 -65
rect 255 -71 259 -67
rect 63 -83 67 -79
<< nsubstratencontact >>
rect 46 14 50 18
rect 57 14 61 18
rect 118 14 122 18
rect 183 14 187 18
rect 234 14 238 18
rect 87 -9 93 -4
rect 150 -9 156 -4
rect 222 -8 229 -3
rect 298 -8 304 -3
rect 98 -68 102 -64
rect 161 -68 166 -63
rect 211 -68 217 -62
rect 286 -68 291 -62
<< labels >>
rlabel metal2 36 -74 36 -74 1 Iref
rlabel metal1 35 16 35 16 1 Vdd
rlabel metal2 45 -68 49 -68 5 Din1
rlabel metal2 107 -68 111 -68 5 Din2
rlabel metal2 175 -68 180 -68 5 Din3
rlabel metal2 243 -68 248 -68 5 Din4
rlabel metal1 311 16 311 16 7 Vdd
rlabel metal1 264 -82 264 -82 1 GND
rlabel metal1 46 -82 46 -82 1 GND
rlabel space 284 -102 284 -93 7 Vout
<< end >>
